//interface definition for 4-bit adder
interface adder_if;
 logic [3:0]a,b;
 logic [4:0] sum;

endinterface